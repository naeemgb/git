
// memory[7] = 32'b000100,00000,00010,00110,00000100010;  // sample
module memoryInstructor (input [31:0]pc,output [31:0]command);
  reg[31:0] memory[0:1023];
  initial begin
		// without any hazard 
		// memory[0] = 32'b10001100000000010000000000000000;  // ld R0 R1 0
		// memory[4] = 32'b10001100000000100000000000000001; // ld R0 R2 1
		// memory[8] = 32'b10001100000000110000000000000010;  // ld R0 R3 2
		// memory[12] = 32'b10001100001001000000000000000010;  // ld R1 R4 2
		// memory[16] = 32'b00000000001000100010100000100000;  // Add R1 R2 R5
		// memory[20] = 32'b00000000011000100011000000100010;  // sub R3 R2 R6
		// memory[24] = 32'b00000000001000100011100000101010;  // slt R1 R2 R7
		// // memory[7] = 32'b00010000000000100011000000100010;  // beg R0 R2 ??		should not jump
		// memory[32] = 32'b00010100000000100000000000000010;  // bne R0 R2 36 			 has to jump
		// memory[28] = 32'b00010000000000100000000000000010;  // bne R0 R2 36 			 should not  jump
		// memory[44] = 32'b11111100000000100011000000100010;  // nop
		// memory[48] = 32'b10101100000001110000000000010010;  // sw R0 R5 17

		// // just forwarding unit 
		// memory[52] = 32'b00000000001000110001000000100010;  // sub R1 R3 R2 ==-15
		// memory[56] = 32'b00000000010001010110000000100100;  // and R2 R5 R12 == -1
		// memory[60] = 32'b00000000110000100110100000100101;  // or R6 R2 R13 == -11
		// memory[64] = 32'b00000000010000100111000000100000;  // add R2 R2 R14 == -30
		// memory[68] = 32'b10101100010011110000000000011000;  // sw R2 R15 24  == mem[9] = R15

		// // hazard unit
		// memory[72] = 32'b10001100001000100000000000010000;  // lw R1 R2 16 == R2 = mem[26] = 59
		// memory[76] = 32'b00000000010001011000000000100000;  // add R2 R5 R16 = 74
		// memory[80] = 32'b00000001100000101000100000100101;  // or R12 R2 R17 = 58

		//***********************************************************************************************************
		//finding maximum number in an array
		// memory[0] = 32'b10001100000000100000001111100111; // load size of array from memory[999]
		// memory[4] = 32'b00000000000000000001100000100000; // set R3 to zero , R3 counts array
		// memory[8] = 32'b00000000000000000010000000100000; // set R4 to zero , R4 holds maximum number 
		// memory[12] = 32'b11111100000000000000000000000000; // nop
		// memory[16] = 32'b00010000010000110000000000001000; // beq if R3 == R2 to end of commands
		// memory[20] = 32'b10001100011001100000001111101000; // load array[R3 + 1000] in R6
		// memory[24] = 32'b00000000100001100010100000101010; // set R5 to 1 if R4 < R6
		// memory[28] = 32'b11111100000000000000000000000000; // nop
		// memory[32] = 32'b11111100000000000000000000000000; // nop
		// memory[36] = 32'b00010000000001010000000000000001; // beq if R5 == R0 to memory[11] 
		// memory[40] = 32'b00000000000001100010000000100000; // assign R6 to R4
		// memory[44] = 32'b00000000011000010001100000100000; // add R3 = R3 + 1
		// memory[48] = 32'b00001000000000000000000000000011; // jump to memory[3]
		// memory[52] = 32'b10101100010001000000000000000001;  // sample 
		//***************************************************************************

		memory[0] = 32'b10001100000000010000000000000000;//
		memory[4] = 32'b10001100000000100000000000000100;
		memory[8] = 32'b10001100000010000000000000001000;
		memory[12] = 32'b00000000000000010000000000100000;
		memory[16] = 32'b00000000001000100001100000101010;  // sample
		memory[20] = 32'b00000000001000100010000000100101;
		memory[24] = 32'b00000000001000100010100000100100;
		memory[28] = 32'b00000000010000010011000000100010;
		memory[32] = 32'b00000000000000010011100000100000;
		memory[36] = 32'b00000000001000100000100000100000;
		memory[40] = 32'b00000000101001110010100000100000;
		memory[44] = 32'b00000000001001110000100000100000;
		memory[48] = 32'b00000000001001110000100000100000;
		memory[52] = 32'b00010001000001011111111111111011;
		memory[56] = 32'b10101100000000010000000000001100;
		memory[60] = 32'b00001011111111111111111111111111;










    // memory[0] = 16'b0000010111110100;
		//  memory[1] = 16'b0000100111110101;
		//  memory[2] = 16'b1000011000000010;
		//  memory[3] = 16'b0000100111110110;
		//  memory[4] = 16'b1000011000000010;
		//  memory[5] = 16'b0000100111110111;
		//  memory[6] = 16'b1000011000000010;
		//  memory[7] = 16'b0000100111111000;
		//  memory[8] = 16'b1000011000000010;
		//  memory[9] = 16'b0000100111111001;
		//  memory[10] = 16'b1000011000000010;
		//  memory[11] = 16'b0000100111111010;
		//  memory[12] = 16'b1000011000000010;
		//  memory[13] = 16'b0000100111111011;
		//  memory[14] = 16'b1000011000000010;
		//  memory[15] = 16'b0000100111111100;
		//  memory[16] = 16'b1000011000000010;
		//  memory[17] = 16'b0000100111111101;
		//  memory[18] = 16'b1000011000000010;
  end

	assign 	command =memory[pc];
endmodule
